module InstructionMemory(rst, PC, clk, 
	ins_25_0, ins_5_0, ins_15_0, ins_15_11, ins_20_16, ins_25_21, ins_31_26, ins_10_6, ins_26);
input rst;
input[31:0] PC;
reg [7:0] data [32767:0];
input clk;
output reg[25:0] ins_25_0;
output reg[5:0] ins_5_0;
output reg[15:0] ins_15_0;
output reg[4:0] ins_15_11;
output reg[4:0] ins_20_16;
output reg[4:0] ins_25_21; 
output reg[5:0] ins_31_26;
output reg[4:0] ins_10_6;
output reg ins_26;
reg[31:0] temp;
reg[7:0] i; 


always @(posedge clk or PC) begin
if (rst) begin
data[0]=8'h8C; data[1]=8'h83; data[2]=8'h00; data[3]=8'h0A;
data[4]=8'h14; data[5]=8'h61; data[6]=8'h00; data[7]=8'h04;
data[8]=8'h20; data[9]=8'h06; data[10]=8'h00; data[11]=8'h02;
data[24]=8'h20; data[25]=8'h05; data[26]=8'h00; data[27]=8'h02;


//data[0]=8'h20; data[1]=8'h01; data[2]=8'h00; data[3]=8'h01;
//data[4]=8'h8C; data[5]=8'h1E; data[6]=8'h00; data[7]=8'h32; 
//data[8]=8'h20; data[9]=8'h02; data[10]=8'h00; data[11]=8'h21;
//data[12]=8'h10; data[13]=8'h22; data[14]=8'h00; data[15]=8'h08;
//data[16]=8'h33; data[17]=8'hC4; data[18]=8'h00; data[19]=8'h01;
//data[20]=8'h14; data[21]=8'h80; data[22]=8'h00; data[23]=8'h02;
//data[24]=8'h21; data[25]=8'h4A; data[26]=8'h00; data[27]=8'h01;
//data[28]=8'h08; data[29]=8'h00; data[30]=8'h00; data[31]=8'h09;
//data[32]=8'h21; data[33]=8'h29; data[34]=8'h00; data[35]=8'h01;
//data[36]=8'h20; data[37]=8'h21; data[38]=8'h00; data[39]=8'h01;
//data[40]=8'h00; data[41]=8'h1E; data[42]=8'hF0; data[43]=8'h42;
//data[44]=8'h08; data[45]=8'h00; data[46]=8'h00; data[47]=8'h03;
//data[48]=8'h90; data[49]=8'h0B; data[50]=8'h00; data[51]=8'h01;

//data[0]=8'h20; data[1]=8'h03; data[2]=8'h00; data[3]=8'h03;
//data[4]=8'h00; data[5]=8'h60; data[6]=8'h20; data[7]=8'h20;
//data[8]=8'h10; data[9]=8'h83; data[10]=8'h00; data[11]=8'h01;
//data[12]=8'h20; data[13]=8'h26; data[14]=8'h00; data[15]=8'h02;
//data[16]=8'h20; data[17]=8'h47; data[18]=8'h00; data[19]=8'h02;

//data[0]=8'h20; data[1]=8'h0F; data[2]=8'h00; data[3]=8'h90;
//data[4]=8'hAC; data[5]=8'h0F; data[6]=8'h00; data[7]=8'h14;
//data[8]=8'h8C; data[9]=8'h08; data[10]=8'h00; data[11]=8'h14;
//data[12]=8'h20; data[13]=8'h09; data[14]=8'h00; data[15]=8'h01;
//data[16]=8'h00; data[17]=8'h00; data[18]=8'h50; data[19]=8'h20;
//data[20]=8'h20; data[21]=8'h0D; data[22]=8'h00; data[23]=8'h01; 
//data[24]=8'h01; data[25]=8'h20; data[26]=8'h58; data[27]=8'h20;
//data[28]=8'h01; data[29]=8'h2A; data[30]=8'h48; data[31]=8'h20;
//data[32]=8'h01; data[33]=8'h60; data[34]=8'h50; data[35]=8'h20;
//data[36]=8'h01; data[37]=8'h28; data[38]=8'h60; data[39]=8'h2A;
//data[40]=8'h11; data[41]=8'h8D; data[42]=8'hFF; data[43]=8'hFB; 
//data[44]=8'h11; data[45]=8'h28; data[46]=8'h00; data[47]=8'h02;
//data[48]=8'h20; data[49]=8'h0D; data[50]=8'h00; data[51]=8'h37;
//data[52]=8'h08; data[53]=8'h00; data[54]=8'h00; data[55]=8'h0F;
//data[56]=8'h20; data[57]=8'h0D; data[58]=8'h00; data[59]=8'h64;
//data[60]=8'hAC; data[61]=8'h0D; data[62]=8'h00; data[63]=8'h18;

//data[0]=8'h90; data[1]=8'h1E; data[2]=8'h00; data[3]=8'h32;
//data[4]=8'h23; data[5]=8'hDE; data[6]=8'h00; data[7]=8'h01;
//data[8]=8'h20; data[9]=8'h01; data[10]=8'h00; data[11]=8'h01;
//data[12]=8'h20; data[13]=8'h06; data[14]=8'h00; data[15]=8'h00;
//data[16]=8'h10; data[17]=8'h3E; data[18]=8'h00; data[19]=8'h0D;
//data[20]=8'h00; data[21]=8'h20; data[22]=8'h10; data[23]=8'h20; 
//data[24]=8'h00; data[25]=8'h20; data[26]=8'h18; data[27]=8'h20;
//data[28]=8'h0C; data[29]=8'h00; data[30]=8'h00; data[31]=8'h0A;
//data[32]=8'h00; data[33]=8'hC4; data[34]=8'h30; data[35]=8'h20;
//data[36]=8'h08; data[37]=8'h00; data[38]=8'h00; data[39]=8'h04;
//data[40]=8'h20; data[41]=8'h04; data[42]=8'h00; data[43]=8'h00; 
//data[44]=8'h20; data[45]=8'h1D; data[46]=8'h00; data[47]=8'h00;
//data[48]=8'h13; data[49]=8'hA3; data[50]=8'h00; data[51]=8'h03;
//data[52]=8'h00; data[53]=8'h82; data[54]=8'h20; data[55]=8'h20;
//data[56]=8'h23; data[57]=8'hBD; data[58]=8'h00; data[59]=8'h01;
//data[60]=8'h08; data[61]=8'h00; data[62]=8'h00; data[63]=8'h0C;
//data[64]=8'h20; data[65]=8'h21; data[66]=8'h00; data[67]=8'h01; 
//data[68]=8'h03; data[69]=8'hE0; data[70]=8'h00; data[71]=8'h08; 
//data[72]=8'h20; data[73]=8'h01; data[74]=8'h00; data[75]=8'h03;
//data[0]=8'h90; data[1]=8'h1E; data[2]=8'h00; data[3]=8'h32;
//data[4]=8'h23; data[5]=8'hDE; data[6]=8'h00; data[7]=8'h01;
//data[8]=8'h20; data[9]=8'h01; data[10]=8'h00; data[11]=8'h01;
//data[12]=8'h20; data[13]=8'h05; data[14]=8'h00; data[15]=8'h00;
//data[16]=8'h10; data[17]=8'h3E; data[18]=8'h00; data[19]=8'h03; 
//data[20]=8'h00; data[21]=8'hA1; data[22]=8'h28; data[23]=8'h20;
//data[24]=8'h20; data[25]=8'h21; data[26]=8'h00; data[27]=8'h01;
//data[28]=8'h08; data[29]=8'h00; data[30]=8'h00; data[31]=8'h04;
//data[32]=8'h20; data[33]=8'h01; data[34]=8'h00; data[35]=8'h01;
//data[36]=8'h20; data[37]=8'h06; data[38]=8'h00; data[39]=8'h00;
//data[40]=8'h10; data[41]=8'h3E; data[42]=8'h00; data[43]=8'h05;
//data[44]=8'h00; data[45]=8'h20; data[46]=8'h10; data[47]=8'h20; 
//data[48]=8'h00; data[49]=8'h20; data[50]=8'h18; data[51]=8'h20;
//data[52]=8'h0C; data[53]=8'h00; data[54]=8'h00; data[55]=8'h6F;
//data[56]=8'h00; data[57]=8'hC4; data[58]=8'h30; data[59]=8'h20;
//data[60]=8'h08; data[61]=8'h00; data[62]=8'h00; data[63]=8'h0A;
//data[64]=8'h20; data[65]=8'h01; data[66]=8'h00; data[67]=8'h03;
//data[68]=8'h20; data[69]=8'h02; data[70]=8'h00; data[71]=8'h01;
//data[72]=8'h20; data[73]=8'h03; data[74]=8'h00; data[75]=8'h01;
//data[76]=8'h10; data[77]=8'h3E; data[78]=8'h00; data[79]=8'h05;
//data[80]=8'h00; data[81]=8'h43; data[82]=8'h20; data[83]=8'h20;
//data[84]=8'h20; data[85]=8'h62; data[86]=8'h00; data[87]=8'h00;
//data[88]=8'h20; data[89]=8'h83; data[90]=8'h00; data[91]=8'h00;
//data[92]=8'h20; data[93]=8'h21; data[94]=8'h00; data[95]=8'h01;
//data[96]=8'h08; data[97]=8'h00; data[98]=8'h00; data[99]=8'h13;
//data[100]=8'h20; data[101]=8'h67; data[102]=8'h00; data[103]=8'h00;
//data[104]=8'h20; data[105]=8'h01; data[106]=8'h00; data[107]=8'h00;
//data[108]=8'h20; data[109]=8'h03; data[110]=8'h00; data[111]=8'h01;
//data[112]=8'h10; data[113]=8'h3E; data[114]=8'h00; data[115]=8'h05;
//data[116]=8'h20; data[117]=8'h22; data[118]=8'h00; data[119]=8'h01; 
//data[120]=8'h0C; data[121]=8'h00; data[122]=8'h00; data[123]=8'h6F;
//data[124]=8'h20; data[125]=8'h83; data[126]=8'h00; data[127]=8'h00;
//data[128]=8'h20; data[129]=8'h21; data[130]=8'h00; data[131]=8'h00;
//data[132]=8'h08; data[133]=8'h00; data[134]=8'h00; data[135]=8'h1C;
//data[136]=8'h20; data[137]=8'h68; data[138]=8'h00; data[139]=8'h00;
//data[140]=8'h20; data[141]=8'h01; data[142]=8'h00; data[143]=8'h01;
//data[144]=8'h8C; data[145]=8'h1E; data[146]=8'h00; data[147]=8'h32; 
//data[148]=8'h20; data[149]=8'h02; data[150]=8'h00; data[151]=8'h21;
//data[152]=8'h10; data[153]=8'h22; data[154]=8'h00; data[155]=8'h08;
//data[156]=8'h33; data[157]=8'hC4; data[158]=8'h00; data[159]=8'h01;
//data[160]=8'h14; data[161]=8'h80; data[162]=8'h00; data[163]=8'h02;
//data[164]=8'h21; data[165]=8'h4A; data[166]=8'h00; data[167]=8'h01;
//data[168]=8'h08; data[169]=8'h00; data[170]=8'h00; data[171]=8'h2C;
//data[172]=8'h21; data[173]=8'h29; data[174]=8'h00; data[175]=8'h01;
//data[176]=8'h20; data[177]=8'h21; data[178]=8'h00; data[179]=8'h01;
//data[180]=8'h00; data[181]=8'h1E; data[182]=8'hF0; data[183]=8'h42;
//data[184]=8'h08; data[185]=8'h00; data[186]=8'h00; data[187]=8'h26;
//data[188]=8'h90; data[189]=8'h0B; data[190]=8'h00; data[191]=8'h01;
//data[192]=8'h90; data[193]=8'h0C; data[194]=8'h00; data[195]=8'h02;
//data[196]=8'h90; data[197]=8'h0D; data[198]=8'h00; data[199]=8'h03;
//data[200]=8'h90; data[201]=8'h0E; data[202]=8'h00; data[203]=8'h04;
//data[204]=8'h90; data[205]=8'h0F; data[206]=8'h00; data[207]=8'h05;
//data[208]=8'h90; data[209]=8'h10; data[210]=8'h00; data[211]=8'h06;
//data[212]=8'h90; data[213]=8'h11; data[214]=8'h00; data[215]=8'h07;
//data[216]=8'h90; data[217]=8'h12; data[218]=8'h00; data[219]=8'h08; 
//data[220]=8'h90; data[221]=8'h13; data[222]=8'h00; data[223]=8'h09;
//data[224]=8'h20; data[225]=8'h01; data[226]=8'h00; data[227]=8'h01;
//data[228]=8'h20; data[229]=8'h04; data[230]=8'h00; data[231]=8'h0A;
//data[232]=8'h10; data[233]=8'h24; data[234]=8'h00; data[235]=8'h2A;
//data[236]=8'h21; data[237]=8'h62; data[238]=8'h00; data[239]=8'h00;
//data[240]=8'h21; data[241]=8'h83; data[242]=8'h00; data[243]=8'h00;
//data[244]=8'h0C; data[245]=8'h00; data[246]=8'h00; data[247]=8'h77; 
//data[248]=8'h20; data[249]=8'h4B; data[250]=8'h00; data[251]=8'h00;
//data[252]=8'h20; data[253]=8'h6C; data[254]=8'h00; data[255]=8'h00;
//data[256]=8'h21; data[257]=8'h82; data[258]=8'h00; data[259]=8'h00;
//data[260]=8'h21; data[261]=8'hA3; data[262]=8'h00; data[263]=8'h00;
//data[264]=8'h0C; data[265]=8'h00; data[266]=8'h00; data[267]=8'h77;
//data[268]=8'h20; data[269]=8'h4C; data[270]=8'h00; data[271]=8'h00;
//data[272]=8'h20; data[273]=8'h6D; data[274]=8'h00; data[275]=8'h00;
//data[276]=8'h21; data[277]=8'hA2; data[278]=8'h00; data[279]=8'h00;
//data[280]=8'h21; data[281]=8'hC3; data[282]=8'h00; data[283]=8'h00;
//data[284]=8'h0C; data[285]=8'h00; data[286]=8'h00; data[287]=8'h77;
//data[288]=8'h20; data[289]=8'h4D; data[290]=8'h00; data[291]=8'h00;
//data[292]=8'h20; data[293]=8'h6E; data[294]=8'h00; data[295]=8'h00;
//data[296]=8'h21; data[297]=8'hC2; data[298]=8'h00; data[299]=8'h00;
//data[300]=8'h21; data[301]=8'hE3; data[302]=8'h00; data[303]=8'h00;
//data[304]=8'h0C; data[305]=8'h00; data[306]=8'h00; data[307]=8'h77;
//data[308]=8'h20; data[309]=8'h4E; data[310]=8'h00; data[311]=8'h00;
//data[312]=8'h20; data[313]=8'h6F; data[314]=8'h00; data[315]=8'h00;
//data[316]=8'h21; data[317]=8'hE2; data[318]=8'h00; data[319]=8'h00; 
//data[320]=8'h22; data[321]=8'h03; data[322]=8'h00; data[323]=8'h00;
//data[324]=8'h0C; data[325]=8'h00; data[326]=8'h00; data[327]=8'h77;
//data[328]=8'h20; data[329]=8'h4F; data[330]=8'h00; data[331]=8'h00;
//data[332]=8'h20; data[333]=8'h70; data[334]=8'h00; data[335]=8'h00;
//data[336]=8'h22; data[337]=8'h02; data[338]=8'h00; data[339]=8'h00;
//data[340]=8'h22; data[341]=8'h23; data[342]=8'h00; data[343]=8'h00;
//data[344]=8'h0C; data[345]=8'h00; data[346]=8'h00; data[347]=8'h77; 
//data[348]=8'h20; data[349]=8'h50; data[350]=8'h00; data[351]=8'h00;
//data[352]=8'h20; data[353]=8'h71; data[354]=8'h00; data[355]=8'h00;
//data[356]=8'h22; data[357]=8'h22; data[358]=8'h00; data[359]=8'h00;
//data[360]=8'h22; data[361]=8'h43; data[362]=8'h00; data[363]=8'h00;
//data[364]=8'h0C; data[365]=8'h00; data[366]=8'h00; data[367]=8'h77;
//data[368]=8'h20; data[369]=8'h51; data[370]=8'h00; data[371]=8'h00;
//data[372]=8'h20; data[373]=8'h72; data[374]=8'h00; data[375]=8'h00;
//data[376]=8'h22; data[377]=8'h42; data[378]=8'h00; data[379]=8'h00;
//data[380]=8'h22; data[381]=8'h63; data[382]=8'h00; data[383]=8'h00;
//data[384]=8'h0C; data[385]=8'h00; data[386]=8'h00; data[387]=8'h77;
//data[388]=8'h20; data[389]=8'h52; data[390]=8'h00; data[391]=8'h00;
//data[392]=8'h20; data[393]=8'h73; data[394]=8'h00; data[395]=8'h00;
//data[396]=8'h20; data[397]=8'h21; data[398]=8'h00; data[399]=8'h01;
//data[400]=8'h08; data[401]=8'h00; data[402]=8'h00; data[403]=8'h3A;
//data[404]=8'h21; data[405]=8'h74; data[406]=8'h00; data[407]=8'h00;
//data[408]=8'h21; data[409]=8'h95; data[410]=8'h00; data[411]=8'h00;
//data[412]=8'h21; data[413]=8'hB6; data[414]=8'h00; data[415]=8'h00;
//data[416]=8'h21; data[417]=8'hD7; data[418]=8'h00; data[419]=8'h00; 
//data[420]=8'h21; data[421]=8'hF8; data[422]=8'h00; data[423]=8'h00;
//data[424]=8'h22; data[425]=8'h19; data[426]=8'h00; data[427]=8'h00;
//data[428]=8'h22; data[429]=8'h3A; data[430]=8'h00; data[431]=8'h00;
//data[432]=8'h22; data[433]=8'h5B; data[434]=8'h00; data[435]=8'h00;
//data[436]=8'h22; data[437]=8'h7C; data[438]=8'h00; data[439]=8'h00;
//data[440]=8'h08; data[441]=8'h00; data[442]=8'h00; data[443]=8'h7D;
//data[444]=8'h20; data[445]=8'h04; data[446]=8'h00; data[447]=8'h00; 
//data[448]=8'h20; data[449]=8'h1D; data[450]=8'h00; data[451]=8'h00;
//data[452]=8'h13; data[453]=8'hA3; data[454]=8'h00; data[455]=8'h03;
//data[456]=8'h00; data[457]=8'h82; data[458]=8'h20; data[459]=8'h20;
//data[460]=8'h23; data[461]=8'hBD; data[462]=8'h00; data[463]=8'h01;
//data[464]=8'h08; data[465]=8'h00; data[466]=8'h00; data[467]=8'h71;
//data[468]=8'h20; data[469]=8'h21; data[470]=8'h00; data[471]=8'h01; 
//data[472]=8'h03; data[473]=8'hE0; data[474]=8'h00; data[475]=8'h08; 
//data[476]=8'h00; data[477]=8'h43; data[478]=8'hF0; data[479]=8'h2A;
//data[480]=8'h17; data[481]=8'hC0; data[482]=8'h00; data[483]=8'h03;
//data[484]=8'h20; data[485]=8'h5D; data[486]=8'h00; data[487]=8'h00;
//data[488]=8'h20; data[489]=8'h62; data[490]=8'h00; data[491]=8'h00;
//data[492]=8'h23; data[493]=8'hA3; data[494]=8'h00; data[495]=8'h00;
//data[496]=8'h03; data[497]=8'hE0; data[498]=8'h00; data[499]=8'h08;
//data[500]=8'h3C; data[501]=8'h01; data[502]=8'hAB; data[503]=8'hCD; 
//data[504]=8'h34; data[505]=8'h22; data[506]=8'h01; data[507]=8'h01;
//data[508]=8'h00; data[509]=8'h22; data[510]=8'h18; data[511]=8'h24;
//data[512]=8'h00; data[513]=8'h22; data[514]=8'h20; data[515]=8'h25;
//data[516]=8'h00; data[517]=8'h22; data[518]=8'hE8; data[519]=8'h27;
//data[520]=8'h28; data[521]=8'h3E; data[522]=8'hFF; data[523]=8'hFF;
//data[524]=8'hA0; data[525]=8'h1E; data[526]=8'h00; data[527]=8'h31;
//data[528]=8'hAC; data[529]=8'h1D; data[530]=8'h00; data[531]=8'h2C;
end
else
begin
		temp = {data[PC[15:0]],data[PC[15:0]+1],data[PC[15:0]+2],data[PC[15:0]+3]};
	end 
end
always @(negedge clk)
begin
ins_25_0 <= temp[25:0];
		ins_5_0 <= temp[5:0];
		ins_15_0 <= temp[15:0];
		ins_15_11 <= temp[15:11];
		ins_20_16 <= temp[20:16];
		ins_25_21 <= temp[25:21]; 
		ins_31_26 <= temp[31:26];
		ins_10_6 <= temp[10:6];
		ins_26 <= temp[26];
end
endmodule
